LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY Final IS 
	PORT
	(
		CLK_BTN :  IN  STD_LOGIC;
		CLK :  IN  STD_LOGIC;
		RESET :  IN  STD_LOGIC;
		DIP1 :  IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
		OUTPUT1 :  OUT  STD_LOGIC;
		OUTPUT2 :  OUT  STD_LOGIC;
		OUTPUT3 :  OUT  STD_LOGIC;
		OUTPUT4 :  OUT  STD_LOGIC;
		sal :  OUT  STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END Final;

ARCHITECTURE bdf_type OF Final IS 

COMPONENT program_counter
	PORT(CLK : IN STD_LOGIC;
		 A_DATA : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 AD : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 OP : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		 OUT_PC : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT extend
	PORT(par2_0 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 par8_6 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 res : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT instruction_memory
	PORT(CLK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;
		 IE : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 I : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT instruction_decoder
	PORT(instruction : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 control_word : OUT STD_LOGIC_VECTOR(19 DOWNTO 0)
	);
END COMPONENT;

COMPONENT unidad_funcional
	PORT(A : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 fs : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		 C : OUT STD_LOGIC;
		 N : OUT STD_LOGIC;
		 Z : OUT STD_LOGIC;
		 F : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT data_memory
	PORT(CLK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;
		 MW : IN STD_LOGIC;
		 Address : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Data_in : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 Data_out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT multiplexer_2_to_1
	PORT(S : IN STD_LOGIC;
		 I0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 I1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 ZERO : OUT STD_LOGIC;
		 Y : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT hexadisplay
	PORT(input_1 : IN STD_LOGIC;
		 dip_1 : IN STD_LOGIC_VECTOR(0 TO 3);
		 dip_2 : IN STD_LOGIC_VECTOR(0 TO 3);
		 dip_3 : IN STD_LOGIC_VECTOR(0 TO 3);
		 dip_4 : IN STD_LOGIC_VECTOR(0 TO 3);
		 output_1 : OUT STD_LOGIC;
		 output_2 : OUT STD_LOGIC;
		 output_3 : OUT STD_LOGIC;
		 output_4 : OUT STD_LOGIC;
		 sal : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END COMPONENT;

COMPONENT register_file
	PORT(CLK : IN STD_LOGIC;
		 RESET : IN STD_LOGIC;
		 RW : IN STD_LOGIC;
		 AA : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 BA : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 D_data_in : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		 DA : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 REG_ADD : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 A_data_out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 B_data_out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		 HEX_OUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT zero_fill
	PORT(z_in : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		 z_out : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END COMPONENT;

COMPONENT branch_control
	PORT(PL : IN STD_LOGIC;
		 JB : IN STD_LOGIC;
		 BC : IN STD_LOGIC;
		 N : IN STD_LOGIC;
		 Z : IN STD_LOGIC;
		 oper : OUT STD_LOGIC_VECTOR(1 DOWNTO 0)
	);
END COMPONENT;

SIGNAL	control_word :  STD_LOGIC_VECTOR(19 DOWNTO 0);
SIGNAL	HEX_OUT :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	I :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_1 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_2 :  STD_LOGIC_VECTOR(1 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_3 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_10 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC_VECTOR(15 DOWNTO 0);
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;


BEGIN 



b2v_inst : program_counter
PORT MAP(CLK => CLK_BTN,
		 A_DATA => SYNTHESIZED_WIRE_15,
		 AD => SYNTHESIZED_WIRE_1,
		 OP => SYNTHESIZED_WIRE_2,
		 OUT_PC => SYNTHESIZED_WIRE_3);


b2v_inst1 : extend
PORT MAP(par2_0 => I(2 DOWNTO 0),
		 par8_6 => I(8 DOWNTO 6),
		 res => SYNTHESIZED_WIRE_1);


b2v_inst10 : instruction_memory
PORT MAP(CLK => CLK_BTN,
		 RESET => RESET,
		 IE => SYNTHESIZED_WIRE_3,
		 I => I);


b2v_inst12 : instruction_decoder
PORT MAP(instruction => I,
		 control_word => control_word);


b2v_inst14 : unidad_funcional
PORT MAP(A => SYNTHESIZED_WIRE_15,
		 B => SYNTHESIZED_WIRE_16,
		 fs => control_word(9 DOWNTO 6),
		 N => SYNTHESIZED_WIRE_13,
		 Z => SYNTHESIZED_WIRE_14,
		 F => SYNTHESIZED_WIRE_10);


b2v_inst15 : data_memory
PORT MAP(CLK => CLK_BTN,
		 RESET => RESET,
		 MW => control_word(3),
		 Address => SYNTHESIZED_WIRE_15,
		 Data_in => SYNTHESIZED_WIRE_16,
		 Data_out => SYNTHESIZED_WIRE_11);


b2v_inst16 : multiplexer_2_to_1
PORT MAP(S => control_word(10),
		 I0 => SYNTHESIZED_WIRE_8,
		 I1 => SYNTHESIZED_WIRE_9,
		 Y => SYNTHESIZED_WIRE_16);


b2v_inst17 : multiplexer_2_to_1
PORT MAP(S => control_word(5),
		 I0 => SYNTHESIZED_WIRE_10,
		 I1 => SYNTHESIZED_WIRE_11,
		 Y => SYNTHESIZED_WIRE_12);


b2v_inst18 : hexadisplay
PORT MAP(input_1 => CLK,
		 dip_1 => HEX_OUT(3 DOWNTO 0),
		 dip_2 => HEX_OUT(7 DOWNTO 4),
		 dip_3 => HEX_OUT(11 DOWNTO 8),
		 dip_4 => HEX_OUT(15 DOWNTO 12),
		 output_1 => OUTPUT1,
		 output_2 => OUTPUT2,
		 output_3 => OUTPUT3,
		 output_4 => OUTPUT4,
		 sal => sal);


b2v_inst19 : register_file
PORT MAP(CLK => CLK_BTN,
		 RESET => RESET,
		 RW => control_word(4),
		 AA => control_word(16 DOWNTO 14),
		 BA => control_word(13 DOWNTO 11),
		 D_data_in => SYNTHESIZED_WIRE_12,
		 DA => control_word(19 DOWNTO 17),
		 REG_ADD => "001",
		 A_data_out => SYNTHESIZED_WIRE_15,
		 B_data_out => SYNTHESIZED_WIRE_8,
		 HEX_OUT => HEX_OUT);


b2v_inst20 : zero_fill
PORT MAP(z_in => I(2 DOWNTO 0),
		 z_out => SYNTHESIZED_WIRE_9);


b2v_inst8 : branch_control
PORT MAP(PL => control_word(2),
		 JB => control_word(1),
		 BC => control_word(0),
		 N => SYNTHESIZED_WIRE_13,
		 Z => SYNTHESIZED_WIRE_14,
		 oper => SYNTHESIZED_WIRE_2);


END bdf_type;