LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY tutorial_altera IS 
	PORT
	(
		A_in :  IN  STD_LOGIC;	
		B_in :  IN  STD_LOGIC;
		C_in :  IN  STD_LOGIC;
		D_in :  IN  STD_LOGIC;
		pin_name1 :  OUT  STD_LOGIC;
		pin_name2 :  OUT  STD_LOGIC;
		pin_name3 :  OUT  STD_LOGIC;
		pin_name9 :  OUT  STD_LOGIC;
		pin_name0 :  OUT  STD_LOGIC;
		pin_name234234 :  OUT  STD_LOGIC;
		fin :  OUT  STD_LOGIC
	);
END tutorial_altera;

ARCHITECTURE bdf_type OF tutorial_altera IS 

SIGNAL	SYNTHESIZED_WIRE_56 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_57 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_58 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_59 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_60 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_61 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_62 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_63 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_26 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_64 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_48 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_51 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_48 <= SYNTHESIZED_WIRE_56 AND C_in;


SYNTHESIZED_WIRE_6 <= SYNTHESIZED_WIRE_56 AND SYNTHESIZED_WIRE_57 AND SYNTHESIZED_WIRE_58;


SYNTHESIZED_WIRE_58 <= NOT(D_in);



SYNTHESIZED_WIRE_7 <= SYNTHESIZED_WIRE_56 AND C_in AND D_in;


pin_name2 <= SYNTHESIZED_WIRE_59 OR SYNTHESIZED_WIRE_6 OR SYNTHESIZED_WIRE_7 OR SYNTHESIZED_WIRE_8;


SYNTHESIZED_WIRE_13 <= SYNTHESIZED_WIRE_56 AND B_in;


SYNTHESIZED_WIRE_12 <= SYNTHESIZED_WIRE_56 AND D_in;


pin_name3 <= SYNTHESIZED_WIRE_60 OR SYNTHESIZED_WIRE_12 OR SYNTHESIZED_WIRE_13 OR SYNTHESIZED_WIRE_59;


SYNTHESIZED_WIRE_62 <= SYNTHESIZED_WIRE_56 AND C_in AND SYNTHESIZED_WIRE_58;


SYNTHESIZED_WIRE_56 <= NOT(A_in);



SYNTHESIZED_WIRE_63 <= SYNTHESIZED_WIRE_56 AND SYNTHESIZED_WIRE_61 AND C_in;


SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_56 AND B_in AND SYNTHESIZED_WIRE_57 AND D_in;


SYNTHESIZED_WIRE_26 <= SYNTHESIZED_WIRE_62 OR SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_60 OR SYNTHESIZED_WIRE_63;


pin_name9 <= SYNTHESIZED_WIRE_59 OR SYNTHESIZED_WIRE_26;


pin_name0 <= SYNTHESIZED_WIRE_60 OR SYNTHESIZED_WIRE_62;


SYNTHESIZED_WIRE_64 <= SYNTHESIZED_WIRE_56 AND B_in AND SYNTHESIZED_WIRE_57;


SYNTHESIZED_WIRE_39 <= SYNTHESIZED_WIRE_56 AND SYNTHESIZED_WIRE_57 AND SYNTHESIZED_WIRE_58;


SYNTHESIZED_WIRE_37 <= SYNTHESIZED_WIRE_56 AND B_in AND SYNTHESIZED_WIRE_58;


pin_name234234 <= SYNTHESIZED_WIRE_64 OR SYNTHESIZED_WIRE_37 OR SYNTHESIZED_WIRE_59 OR SYNTHESIZED_WIRE_39;


fin <= SYNTHESIZED_WIRE_62 OR SYNTHESIZED_WIRE_64 OR SYNTHESIZED_WIRE_59 OR SYNTHESIZED_WIRE_63;


SYNTHESIZED_WIRE_51 <= SYNTHESIZED_WIRE_56 AND B_in AND D_in;


SYNTHESIZED_WIRE_60 <= SYNTHESIZED_WIRE_61 AND SYNTHESIZED_WIRE_57 AND SYNTHESIZED_WIRE_58;


SYNTHESIZED_WIRE_57 <= NOT(C_in);



SYNTHESIZED_WIRE_61 <= NOT(B_in);



pin_name1 <= SYNTHESIZED_WIRE_48 OR SYNTHESIZED_WIRE_60 OR SYNTHESIZED_WIRE_59 OR SYNTHESIZED_WIRE_51;


SYNTHESIZED_WIRE_8 <= SYNTHESIZED_WIRE_56 AND SYNTHESIZED_WIRE_61;


SYNTHESIZED_WIRE_59 <= A_in AND SYNTHESIZED_WIRE_61 AND SYNTHESIZED_WIRE_57;


END bdf_type;